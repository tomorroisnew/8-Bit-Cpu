module Uart()